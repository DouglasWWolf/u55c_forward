/*
================================================================================================
  Vers     Date    Who  Changes
------- ----------------------------------------------------------------------------------------
 1.0.0  21-Jan-26  DWW  Initial creation
================================================================================================
*/

localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 0;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 0;


localparam RTL_TYPE      = 12126;
localparam RTL_SUBTYPE   = 0;
